`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    18:35:36 11/24/2015 
// Design Name: 
// Module Name:    divisor_black 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module divisor_black(
	input wire [1183:0]buffer_envio,
	output reg [7:0]o1,
	output reg [7:0]o2,
	output reg [7:0]o3,
	output reg [7:0]o4,
	output reg [7:0]o5,
	output reg [7:0]o6,
	output reg [7:0]o7,
	output reg [7:0]o8,
	output reg [7:0]o9,
	output reg [7:0]o10,
	output reg [7:0]o11,
	output reg [7:0]o12,
	output reg [7:0]o13,
	output reg [7:0]o14,
	output reg [7:0]o15,
	output reg [7:0]o16,
	output reg [7:0]o17,
	output reg [7:0]o18,
	output reg [7:0]o19,
	output reg [7:0]o20,
	output reg [7:0]o21,
	output reg [7:0]o22,
	output reg [7:0]o23,
	output reg [7:0]o24,
	output reg [7:0]o25,
	output reg [7:0]o26,
	output reg [7:0]o27,
	output reg [7:0]o28,
	output reg [7:0]o29,
	output reg [7:0]o30,
	output reg [7:0]o31,
	output reg [7:0]o32,
	output reg [7:0]o33,
	output reg [7:0]o34,
	output reg [7:0]o35,
	output reg [7:0]o36,
	output reg [7:0]o37,
	output reg [7:0]o38,
	output reg [7:0]o39,
	output reg [7:0]o40,
	output reg [7:0]o41,
	output reg [7:0]o42,
	output reg [7:0]o43,
	output reg [7:0]o44,
	output reg [7:0]o45,
	output reg [7:0]o46,
	output reg [7:0]o47,
	output reg [7:0]o48,
	output reg [7:0]o49,
	output reg [7:0]o50,
	output reg [7:0]o51,
	output reg [7:0]o52,
	output reg [7:0]o53,
	output reg [7:0]o54,
	output reg [7:0]o55,
	output reg [7:0]o56,
	output reg [7:0]o57,
	output reg [7:0]o58,
	output reg [7:0]o59,
	output reg [7:0]o60,
	output reg [7:0]o61,
	output reg [7:0]o62,
	output reg [7:0]o63,
	output reg [7:0]o64,
	output reg [7:0]o65,
	output reg [7:0]o66,
	output reg [7:0]o67,
	output reg [7:0]o68,
	output reg [7:0]o69,
	output reg [7:0]o70,
	output reg [7:0]o71,
	output reg [7:0]o72,
	output reg [7:0]o73,
	output reg [7:0]o74,
	output reg [7:0]o75,
	output reg [7:0]o76,
	output reg [7:0]o77,
	output reg [7:0]o78,
	output reg [7:0]o79,
	output reg [7:0]o80,
	output reg [7:0]o81,
	output reg [7:0]o82,
	output reg [7:0]o83,
	output reg [7:0]o84,
	output reg [7:0]o85,
	output reg [7:0]o86,
	output reg [7:0]o87,
	output reg [7:0]o88,
	output reg [7:0]o89,
	output reg [7:0]o90,
	output reg [7:0]o91,
	output reg [7:0]o92,
	output reg [7:0]o93,
	output reg [7:0]o94,
	output reg [7:0]o95,
	output reg [7:0]o96,
	output reg [7:0]o97,
	output reg [7:0]o98,
	output reg [7:0]o99,
	output reg [7:0]o100,
	output reg [7:0]o101,
	output reg [7:0]o102,
	output reg [7:0]o103,
	output reg [7:0]o104,
	output reg [7:0]o105,
	output reg [7:0]o106,
	output reg [7:0]o107,
	output reg [7:0]o108,
	output reg [7:0]o109,
	output reg [7:0]o110,
	output reg [7:0]o111,
	output reg [7:0]o112,
	output reg [7:0]o113,
	output reg [7:0]o114,
	output reg [7:0]o115,
	output reg [7:0]o116,
	output reg [7:0]o117,
	output reg [7:0]o118,
	output reg [7:0]o119,
	output reg [7:0]o120,
	output reg [7:0]o121,
	output reg [7:0]o122,
	output reg [7:0]o123,
	output reg [7:0]o124,
	output reg [7:0]o125,
	output reg [7:0]o126,
	output reg [7:0]o127,
	output reg [7:0]o128,
	output reg [7:0]o129,
	output reg [7:0]o130,
	output reg [7:0]o131,
	output reg [7:0]o132,
	output reg [7:0]o133,
	output reg [7:0]o134,
	output reg [7:0]o135,
	output reg [7:0]o136,
	output reg [7:0]o137,
	output reg [7:0]o138,
	output reg [7:0]o139,
	output reg [7:0]o140,
	output reg [7:0]o141,
	output reg [7:0]o142,
	output reg [7:0]o143,
	output reg [7:0]o144,
	output reg [7:0]o145,
	output reg [7:0]o146,
	output reg [7:0]o147,
	output reg [7:0]o148
 );

always@(*)
begin
	o1 <= buffer_envio[7:0];
	o2 <= buffer_envio[15:8];
	o3 <= buffer_envio[23:16];
	o4 <= buffer_envio[31:24];
	o5 <= buffer_envio[39:32];
	o6 <= buffer_envio[47:40];
	o7 <= buffer_envio[55:48];
	o8 <= buffer_envio[63:56];
	o9 <= buffer_envio[71:64];
	o10 <= buffer_envio[79:72];
	o11 <= buffer_envio[87:80];
	o12 <= buffer_envio[95:88];
	o13 <= buffer_envio[103:96];
	o14 <= buffer_envio[111:104];
	o15 <= buffer_envio[119:112];
	o16 <= buffer_envio[127:120];
	o17 <= buffer_envio[135:128];
	o18 <= buffer_envio[143:136];
	o19 <= buffer_envio[151:144];
	o20 <= buffer_envio[159:152];
	o21 <= buffer_envio[167:160];
	o22 <= buffer_envio[175:168];
	o23 <= buffer_envio[183:176];
	o24 <= buffer_envio[191:184];
	o25 <= buffer_envio[199:192];
	o26 <= buffer_envio[207:200];
	o27 <= buffer_envio[215:208];
	o28 <= buffer_envio[223:216];
	o29 <= buffer_envio[231:224];
	o30 <= buffer_envio[239:232];
	o31 <= buffer_envio[247:240];
	o32 <= buffer_envio[255:248];
	o33 <= buffer_envio[263:256];
	o34 <= buffer_envio[271:264];
	o35 <= buffer_envio[279:272];
	o36 <= buffer_envio[287:280];
	o37 <= buffer_envio[295:288];
	o38 <= buffer_envio[303:296];
	o39 <= buffer_envio[311:304];
	o40 <= buffer_envio[319:312];
	o41 <= buffer_envio[327:320];
	o42 <= buffer_envio[335:328];
	o43 <= buffer_envio[343:336];
	o44 <= buffer_envio[351:344];
	o45 <= buffer_envio[359:352];
	o46 <= buffer_envio[367:360];
	o47 <= buffer_envio[375:368];
	o48 <= buffer_envio[383:376];
	o49 <= buffer_envio[391:384];
	o50 <= buffer_envio[399:392];
	o51 <= buffer_envio[407:400];
	o52 <= buffer_envio[415:408];
	o53 <= buffer_envio[423:416];
	o54 <= buffer_envio[431:424];
	o55 <= buffer_envio[439:432];
	o56 <= buffer_envio[447:440];
	o57 <= buffer_envio[455:448];
	o58 <= buffer_envio[463:456];
	o59 <= buffer_envio[471:464];
	o60 <= buffer_envio[479:472];
	o61 <= buffer_envio[487:480];
	o62 <= buffer_envio[495:488];
	o63 <= buffer_envio[503:496];
	o64 <= buffer_envio[511:504];
	o65 <= buffer_envio[519:512];
	o66 <= buffer_envio[527:520];
	o67 <= buffer_envio[535:528];
	o68 <= buffer_envio[543:536];
	o69 <= buffer_envio[551:544];
	o70 <= buffer_envio[559:552];
	o71 <= buffer_envio[567:560];
	o72 <= buffer_envio[575:568];
	o73 <= buffer_envio[583:576];
	o74 <= buffer_envio[591:584];
	o75 <= buffer_envio[599:592];
	o76 <= buffer_envio[607:600];
	o77 <= buffer_envio[615:608];
	o78 <= buffer_envio[623:616];
	o79 <= buffer_envio[631:624];
	o80 <= buffer_envio[639:632];
	o81 <= buffer_envio[647:640];
	o82 <= buffer_envio[655:648];
	o83 <= buffer_envio[663:656];
	o84 <= buffer_envio[671:664];
	o85 <= buffer_envio[679:672];
	o86 <= buffer_envio[687:680];
	o87 <= buffer_envio[695:688];
	o88 <= buffer_envio[703:696];
	o89 <= buffer_envio[711:704];
	o90 <= buffer_envio[719:712];
	o91 <= buffer_envio[727:720];
	o92 <= buffer_envio[735:728];
	o93 <= buffer_envio[743:736];
	o94 <= buffer_envio[751:744];
	o95 <= buffer_envio[759:752];
	o96 <= buffer_envio[767:760];
	o97 <= buffer_envio[775:768];
	o98 <= buffer_envio[783:776];
	o99 <= buffer_envio[791:784];
	o100 <= buffer_envio[799:792];
	o101 <= buffer_envio[807:800];
	o102 <= buffer_envio[815:808];
	o103 <= buffer_envio[823:816];
	o104 <= buffer_envio[831:824];
	o105 <= buffer_envio[839:832];
	o106 <= buffer_envio[847:840];
	o107 <= buffer_envio[855:848];
	o108 <= buffer_envio[863:856];
	o109 <= buffer_envio[871:864];
	o110 <= buffer_envio[879:872];
	o111 <= buffer_envio[887:880];
	o112 <= buffer_envio[895:888];
	o113 <= buffer_envio[903:896];
	o114 <= buffer_envio[911:904];
	o115 <= buffer_envio[919:912];
	o116 <= buffer_envio[927:920];
	o117 <= buffer_envio[935:928];
	o118 <= buffer_envio[943:936];
	o119 <= buffer_envio[951:944];
	o120 <= buffer_envio[959:952];
	o121 <= buffer_envio[967:960];
	o122 <= buffer_envio[975:968];
	o123 <= buffer_envio[983:976];
	o124 <= buffer_envio[991:984];
	o125 <= buffer_envio[999:992];
	o126 <= buffer_envio[1007:1000];
	o127 <= buffer_envio[1015:1008];
	o128 <= buffer_envio[1023:1016];
	o129 <= buffer_envio[1031:1024];
	o130 <= buffer_envio[1039:1032];
	o131 <= buffer_envio[1047:1040];
	o132 <= buffer_envio[1055:1048];
	o133 <= buffer_envio[1063:1056];
	o134 <= buffer_envio[1071:1064];
	o135 <= buffer_envio[1079:1072];
	o136 <= buffer_envio[1087:1080];
	o137 <= buffer_envio[1095:1088];
	o138 <= buffer_envio[1103:1096];
	o139 <= buffer_envio[1111:1104];
	o140 <= buffer_envio[1119:1112];
	o141 <= buffer_envio[1127:1120];
	o142 <= buffer_envio[1135:1128];
	o143 <= buffer_envio[1143:1136];
	o144 <= buffer_envio[1151:1144];
	o145 <= buffer_envio[1159:1152];
	o146 <= buffer_envio[1167:1160];
	o147 <= buffer_envio[1175:1168];
	o148 <= buffer_envio[1183:1176];
end

endmodule
