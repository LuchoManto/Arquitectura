`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    19:45:18 08/24/2015 
// Design Name: 
// Module Name:    pruebacarga 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module pruebacarga(
	input wire [7:0]i_bit,
	output wire [7:0]o_led
    );
	 
	 assign o_led = i_bit;
	 

endmodule
