`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    10:18:19 09/18/2015 
// Design Name: 
// Module Name:    ejercicio_11 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module ejercicio_11(
	input wire i_signal;
	output reg o_periodo;
	
	input wire clk;
    );
	 
	 reg cuenta;
	 
	 
	 always@(posedge clock)
	 begin
	 
	 if(posedge i_signal)
	 begin
	 
	 
	 end
	 
	 end


endmodule
